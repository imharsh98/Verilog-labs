/********************************************************************************************
Copyright 2019 - Maven Silicon Softech Pvt Ltd. 
 
All Rights Reserved.

This source code is an unpublished work belongs to Maven Silicon Softech Pvt Ltd.

It is not to be shared with or used by any third parties who have not enrolled for our paid training 

courses or received any written authorization from Maven Silicon.


Webpage     :      www.maven-silicon.com

Filename    :	   mux4_1_tb.v   

Description :      Mux 4:1 Testbench

Author Name :      Susmita

Version     :      1.0
*********************************************************************************************/

module mux4_1_tb();

   //Step1 : Write down the variables required for testbench		
								
   //Step2 : Instantiate the Design 

   //Step3 : Declare a task to initialize inputs of DUT to 0 

   //Step4 : Declare  tasks with arguments for driving stimulus to DUT 

   //Step5 : Call the tasks from procedural process 

   //Step6 : Use $monitor task to display inputs and outputs

   //Step7 : Use $finish task to terminate the simulation at 100ns

   
endmodule

